library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

use work.core_pkg.all;
use work.op_pkg.all;

entity ctrl is
	port (
		clk         : in std_logic;
		res_n       : in std_logic;
		stall       : in std_logic;

		stall_fetch : out std_logic;
		stall_dec   : out std_logic;
		stall_exec  : out std_logic;
		stall_mem   : out std_logic;
		stall_wb    : out std_logic;

		flush_fetch : out std_logic;
		flush_dec   : out std_logic;
		flush_exec  : out std_logic;
		flush_mem   : out std_logic;
		flush_wb    : out std_logic;

		-- from FWD
		wb_op_exec  : in  wb_op_type;
		exec_op_dec : in  exec_op_type;

		pcsrc_in : in std_logic;
		pcsrc_out : out std_logic
	);
end entity;

architecture rtl of ctrl is
	signal load_hazard : std_logic := '0';
begin
	load_hazard <= '1' when wb_op_exec.write = '1' and wb_op_exec.src = WBS_MEM and
				(wb_op_exec.rd = exec_op_dec.rs1 or wb_op_exec.rd = exec_op_dec.rs2) 
			else '0';

	flush_wb    <= '0'; 

	flush_fetch <= pcsrc_in; 
	flush_dec   <= pcsrc_in;
	flush_exec  <= pcsrc_in or load_hazard;
	flush_mem   <= pcsrc_in;   

	stall_fetch <= stall or load_hazard;
	stall_dec   <= stall or load_hazard;
	stall_exec  <= stall;
	stall_mem   <= stall;
	stall_wb    <= stall;
	
	pcsrc_out <= pcsrc_in;

end architecture;
